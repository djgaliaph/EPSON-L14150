��[ G r o u p T i t l e ]  
 P r i n t e r D r i v e r G r o u p 	 	 = " S k r i v a r d r i v r u t i n e r   o c h   - v e r k t y g "  
 S c a n n e r G r o u p 	 	 	 = " S k a n n e r d r i v r u t i n "  
 S c a n n e r U t i l i t y G r o u p 	 	 = " S k a n n e r v e r k t y g "  
 F a x G r o u p 	 	 	 = " F a x v e r k t y g "  
 M a n u a l G r o u p 	 	 	 = " H a n d b � c k e r "  
 U t i l i t y G r o u p 	 	 	 = " S u p p o r t v e r k t y g "  
 P h o t o P l u s G r o u p 	 	 	 = " E p s o n   P h o t o + "  
 S c a n S m a r t G r o u p 	 	 	 = " E p s o n   S c a n S m a r t "  
 S o f t w a r e U p d a t e r G r o u p 	 	 = " S o f t w a r e   U p d a t e r "  
 P L o g G r o u p 	 	 	 = " E p s o n   C u s t o m e r   R e s e a c h "  
 S t a t u s M o n i t o r G r o u p 	 	 = " S t a t u s   M o n i t o r "  
 D o c C a p G r o u p 	 	 	 = " D o c u m e n t   C a p t u r e   P r o "  
 D o c C a p G r o u p _ m 	 	 	 = " D o c u m e n t   C a p t u r e "  
 C l o u d G r o u p 	 	 	 = " C l o u d   S o f t w a r e "  
 P S G r o u p 	 	 	 	 = " P S   ( P o s t S c r i p t )   D r i c e r "  
 N e t w a r e G r o u p 	 	 	 = " A d m i n i s t r a t � r s p r o g r a m "  
  
 [ G r o u p D e s c r i p t i o n ]  
 P r i n t e r D r i v e r G r o u p 	 	 = " "  
 S c a n n e r G r o u p 	 	 	 = " "  
 S c a n n e r U t i l i t y G r o u p 	 	 = " "  
 F a x G r o u p 	 	 	 = " "  
 M a n u a l G r o u p 	 	 	 = " "  
 U t i l i t y G r o u p 	 	 	 = " "  
 P h o t o P l u s G r o u p 	 	 	 = " "  
 S c a n S m a r t G r o u p 	 	 	 = " "  
 S o f t w a r e U p d a t e r G r o u p 	 	 = " "  
 P L o g G r o u p 	 	 	 = " "  
 S t a t u s M o n i t o r G r o u p 	 	 = " "  
 D o c C a p G r o u p 	 	 	 = " "  
 C l o u d G r o u p 	 	 	 = " "  
 P S G r o u p 	 	 	 	 = " "  
 N e t w a r e G r o u p 	 	 	 = " "  
  
 [ S o f t w a r e N a m e ]  
 P r i n t e r D r i v e r x 6 4   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 6 4 _ L P   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 _ L P   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r   	 	 = " S k r i v a r d r i v r u t i n "  
 S c a n n e r D r i v e r   	 	 = " S k a n n e r d r i v r u t i n "  
 E p s o n S c a n O C R C o m p o n e n t   	 = " E p s o n   S c a n   2   O C R   C o m p o n e n t "  
 E p s o n S c a n P D F E x t e n s i o n s   	 = " E p s o n   S c a n   2   P D F   E x t e n s i o n s "  
 E v e n t M a n a g e r   	 	 = " E v e n t   M a n a g e r "  
 D o c u m e n t C a p t u r e   	 = " D o c u m e n t   C a p t u r e   P r o "  
 D o c u m e n t C a p t u r e P r o V 2   	 = " D o c u m e n t   C a p t u r e   P r o "  
 M y E P S O N P o r t a l   	 	 = " M y E P S O N   P o r t a l "  
 D o w n l o a d N a v i g a t o r   	 = " S o f t w a r e   U p d a t e r "  
 E p s o n N e t P r i n t   	 	 = " E p s o n N e t   P r i n t "  
 E p s o n N e t S e t u p 	 	 = " E p s o n N e t   S e t u p "  
 E p s o n N e t C o n f i g   	 	 = " E p s o n N e t   C o n f i g "  
 M a n u a l P a c k a g e   	 	 = " M a n u e l l t "  
 M a n u a l L a u n c h e r   	 	 = " S t a r t p r o g r a m   f � r   h a n d b o k "  
 M a n u a l D a t a   	 	 = " M a n u e l l t "  
 M a n u a l D a t a S c n   	 	 = " M a n u e l l t "  
 E p s o n C o n n e c t S h o r t c u t   	 = " E p s o n   C o n n e c t   S i t e "  
 F a x U t i l i t y   	 	 = " F a x   U t i l i t y "  
 F a x U t i l i t y W   	 	 = " F a x   U t i l i t y "  
 P h o t o P l u s   	 	 = " E p s o n   P h o t o + "  
 P h o t o P l u s X V   	 	 = " E p s o n   P h o t o + "  
 S c a n S m a r t   	 	 = " E p s o n   S c a n S m a r t "  
 S c a n S m a r t W R   	 	 = " E p s o n   S c a n S m a r t "  
 S u p p o r t L i n k   	 	 = " L � n k   t i l l   A n v � n d a r h a n d b o k "  
 F a s t F o t o   	 	 = " F a s t F o t o "  
 F a s t F o t o 2   	 	 = " F a s t F o t o "  
 S t a t u s M o n i t o r x 6 4 	 = " S t a t u s   M o n i t o r "  
 S t a t u s M o n i t o r x 8 6 	 = " S t a t u s   M o n i t o r "  
 S t a t u s M o n i t o r 3 	 	 = " S t a t u s   M o n i t o r "  
 C o n n e c t C h e c k e r   	 	 = " E p s o n   C o n n e c t i o n   C h e c k e r "  
 F A X 1   	 	 	 = " F a x   U t i l i t y "  
 I C A 1   	 	 	 = " I C A   D r i v e r "  
 D C 1   	 	 	 = " D o c u m e n t   C a p t u r e "  
 M A N U A L 1   	 	 = " S t a r t p r o g r a m   f � r   h a n d b o k "  
 E P S O N   S o f t w a r e   U p d a t e r 2   = " S o f t w a r e   U p d a t e r "  
 S c a n S m a r t I J P 	 	 	 = " E p s o n   S c a n S m a r t "  
 D o c u m e n t C a p t u r e P r o V 2 I J P 	 	 = " D o c u m e n t   C a p t u r e   P r o "  
 P r i n t e r D r i v e r x 6 4 _ L a b e l   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 _ L a b e l   	 = " S k r i v a r d r i v r u t i n "  
  
 [ S o f t w a r e N a m e _ a r t i c l e ]  
 P r i n t e r D r i v e r x 6 4   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 6 4 _ L P   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 _ L P   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r   	 	 = " S k r i v a r d r i v r u t i n "  
 S c a n n e r D r i v e r   	 	 = " S k a n n e r d r i v r u t i n "  
 E p s o n S c a n O C R C o m p o n e n t   	 = " E p s o n   S c a n   2   O C R   C o m p o n e n t "  
 E p s o n S c a n P D F E x t e n s i o n s   	 = " E p s o n   S c a n   2   P D F   E x t e n s i o n s "  
 E v e n t M a n a g e r   	 	 = " E v e n t   M a n a g e r "  
 D o c u m e n t C a p t u r e   	 = " D o c u m e n t   C a p t u r e   P r o "  
 D o c u m e n t C a p t u r e P r o V 2   	 = " D o c u m e n t   C a p t u r e   P r o "  
 M y E P S O N P o r t a l   	 	 = " M y E P S O N   P o r t a l "  
 D o w n l o a d N a v i g a t o r   	 = " S o f t w a r e   U p d a t e r "  
 E p s o n N e t P r i n t   	 	 = " E p s o n N e t   P r i n t "  
 E p s o n N e t S e t u p 	 	 = " E p s o n N e t   S e t u p "  
 E p s o n N e t C o n f i g   	 	 = " E p s o n N e t   C o n f i g "  
 M a n u a l P a c k a g e   	 	 = " M a n u e l l t "  
 M a n u a l L a u n c h e r   	 	 = " S t a r t p r o g r a m   f � r   h a n d b o k "  
 M a n u a l D a t a   	 	 = " M a n u e l l t "  
 M a n u a l D a t a S c n   	 	 = " M a n u e l l t "  
 E p s o n C o n n e c t S h o r t c u t   	 = " E p s o n   C o n n e c t   S i t e "  
 F a x U t i l i t y   	 	 = " F a x   U t i l i t y "  
 F a x U t i l i t y W   	 	 = " F a x   U t i l i t y "  
 P h o t o P l u s   	 	 = " E p s o n   P h o t o + "  
 P h o t o P l u s X V   	 	 = " E p s o n   P h o t o + "  
 S c a n S m a r t   	 	 = " E p s o n   S c a n S m a r t "  
 S c a n S m a r t W R   	 	 = " E p s o n   S c a n S m a r t "  
 S u p p o r t L i n k   	 	 = " L � n k   t i l l   A n v � n d a r h a n d b o k "  
 F a s t F o t o   	 	 = " F a s t F o t o "  
 F a s t F o t o 2   	 	 = " F a s t F o t o "  
 S t a t u s M o n i t o r x 6 4 	 = " S t a t u s   M o n i t o r "  
 S t a t u s M o n i t o r x 8 6 	 = " S t a t u s   M o n i t o r "  
 S t a t u s M o n i t o r 3 	 	 = " S t a t u s   M o n i t o r "  
 C o n n e c t C h e c k e r   	 	 = " E p s o n   C o n n e c t i o n   C h e c k e r "  
 F A X 1   	 	 	 = " F a x   U t i l i t y "  
 I C A 1   	 	 	 = " I C A   D r i v e r "  
 D C 1   	 	 	 = " D o c u m e n t   C a p t u r e "  
 M A N U A L 1   	 	 = " S t a r t p r o g r a m   f � r   h a n d b o k "  
 E P S O N   S o f t w a r e   U p d a t e r 2   = " S o f t w a r e   U p d a t e r "  
 S c a n S m a r t I J P 	 	 	 = " E p s o n   S c a n S m a r t "  
 D o c u m e n t C a p t u r e P r o V 2 I J P 	 	 = " D o c u m e n t   C a p t u r e   P r o "  
 P r i n t e r D r i v e r x 6 4 _ L a b e l   	 = " S k r i v a r d r i v r u t i n "  
 P r i n t e r D r i v e r x 8 6 _ L a b e l   	 = " S k r i v a r d r i v r u t i n "  
  
 [ S o f t w a r e D e s c r i p t i o n ]  
 P r i n t e r D r i v e r x 6 4   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 P r i n t e r D r i v e r x 8 6   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 P r i n t e r D r i v e r x 6 4 _ L P   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 P r i n t e r D r i v e r x 8 6 _ L P   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 P r i n t e r D r i v e r   	 	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 S c a n n e r D r i v e r   	 	 = " D e t   l � t e r   d i g   k o n t r o l l e r a   a l l a   a s p e k t e r   a v   s k a n n i n g ,   s k a n n i n g s l � g e ,   f � r g ,   u p p l � s n i n g ,   f o r m a t   a t t   s p a r a   i   o c h   s �   v i d a r e .   ( P r o g r a m v a r u k r a v ) "  
 E p s o n S c a n O C R C o m p o n e n t   	 = " D e t t a   t i l l � g g s p r o g r a m   s p a r a r   s k a n n a d e   b i l d e r   s o m   s � k b a r a   P D F - f i l e r . "  
 E p s o n S c a n P D F E x t e n s i o n s   	 = " D e t t a   t i l l � g g s p r o g r a m   l � s e n o r d s k y d d a r   e n   s k a n n a d   b i l d   s o m   s p a r a s   i   P D F - f o r m a t . "  
 E v e n t M a n a g e r   	 	 = " D e t   l � t e r   d i g   a n v � n d a   s k a n n i n g   f r � n   p r o d u k t e n s   k o n t r o l l p a n e l . "  
 D o c u m e n t C a p t u r e   	 = " D e t   l � t e r   d i g   h a n t e r a   s k a n n a d e   d o k u m e n t   o c h   s p a r a   d e m   s o m   f i l e r   f � r   a t t   s e d a n   s k i c k a   d e m   t i l l   F T P ,   e n   s k r i v a r e   e l l e r   m o l n e t . "  
 D o c u m e n t C a p t u r e P r o V 2   	 = " D e t   l � t e r   d i g   h a n t e r a   s k a n n a d e   d o k u m e n t   o c h   s p a r a   d e m   s o m   f i l e r   f � r   a t t   s e d a n   s k i c k a   d e m   t i l l   F T P ,   e n   s k r i v a r e   e l l e r   m o l n e t . "  
 M y E P S O N P o r t a l   	 	 = " D e t   l � t e r   d i g   f e l s � k a   u t s k r i f t s p r o b l e m   o c h   d e t   s k i c k a r   d i g   s t u n d t a l s   u p p d a t e r i n g a r   s o m   e x e m p e l v i s   s � r s k i l d a   k a m p a n j e r   f r � n   E p s o n . "  
 D o w n l o a d N a v i g a t o r   	 = " D e t   l � t e r   d i g   u p p d a t e r a   d i n   p r o d u k t s   p r o g r a m v a r a   t i l l   d e n   s e n a s t e   v e r s i o n e n . "  
 E P S O N   S o f t w a r e   U p d a t e r 2   = " D e t   l � t e r   d i g   u p p d a t e r a   d i n   p r o d u k t s   p r o g r a m v a r a   t i l l   d e n   s e n a s t e   v e r s i o n e n . "  
 E p s o n N e t P r i n t   	 	 = " E p s o n N e t   P r i n t "  
 E p s o n N e t S e t u p 	 	 = " E p s o n N e t   S e t u p "  
 E p s o n N e t C o n f i g   	 	 = " D e t   l � t e r   a d m i n i s t r a t � r e r   k o n f i g u r e r a   n � t v e r k s g r � n s s n i t t s i n s t � l l n i n g a r   s o m   T C P / I P   o c h   s �   v i d a r e . "  
 M a n u a l P a c k a g e   	 	 = " D e n   b e r � t t a r   h u r   d u   a n v � n d e r ,   u n d e r h � l l e r   o c h   f e l s � k e r   d i n   p r o d u k t . "  
 M a n u a l L a u n c h e r   	 	 = " D e t   s t a r t a r   E p s o n - b r u k s a n v i s n i n g a r   p �   d i n   d a t o r ,   f r � n   E p s o n - w e b b p l a t s e n . "  
 M a n u a l D a t a   	 	 = " D e n   b e r � t t a r   h u r   d u   a n v � n d e r ,   u n d e r h � l l e r   o c h   f e l s � k e r   d i n   p r o d u k t . "  
 M a n u a l D a t a S c n   	 	 = " D e n   b e r � t t a r   h u r   d u   a n v � n d e r ,   u n d e r h � l l e r   o c h   f e l s � k e r   d i n   p r o d u k t . "  
 F a x U t i l i t y   	 	 = " D e t   l � t e r   d i g   s k i c k a   f a x   f r � n   d i n   d a t o r   e l l e r   h a n t e r a   e n   t e l e f o n b o k . "  
 F a x U t i l i t y W   	 	 = " D e t   l � t e r   d i g   s k i c k a   f a x   f r � n   d i n   d a t o r   e l l e r   h a n t e r a   e n   t e l e f o n b o k . "  
 F A X 1   	 	 	 = " D e t   l � t e r   d i g   s k i c k a   f a x   f r � n   d i n   d a t o r   e l l e r   h a n t e r a   e n   t e l e f o n b o k . "  
 P h o t o P l u s   	 	 = " D e n   l � t e r   d i g   s k r i v a   u t   f o t o n   e n k e l t ,   m e d   e t t   u r v a l   a v   m a l l a r ,   o c h   d e t   g � r   o c k s �   a t t   l � g g a   t i l l   b o k s t � v e r   o c h   s t � m p l a r . "  
 P h o t o P l u s X V   	 	 = " D e n   l � t e r   d i g   s k r i v a   u t   f o t o n   e n k e l t ,   m e d   e t t   u r v a l   a v   m a l l a r ,   o c h   d e t   g � r   o c k s �   a t t   l � g g a   t i l l   b o k s t � v e r   o c h   s t � m p l a r . "  
 S c a n S m a r t   	 	 = " D e t   l � t e r   d i g   s k a n n a   d e t   u r s p r u n g l i g a   d o k u m e n t e t   o c h   s e d a n   f � l j a   i n s t r u k t i o n e r n a   p �   s k � r m e n   f � r   a t t   s p a r a   e l l e r   s k i c k a   d e n   s k a n n a d e   b i l d e n . "  
 S c a n S m a r t W R   	 	 = " D e t   l � t e r   d i g   s k a n n a   d e t   u r s p r u n g l i g a   d o k u m e n t e t   o c h   s e d a n   f � l j a   i n s t r u k t i o n e r n a   p �   s k � r m e n   f � r   a t t   s p a r a   e l l e r   s k i c k a   d e n   s k a n n a d e   b i l d e n . "  
 S u p p o r t L i n k   	 	 = " D e n   b e r � t t a r   h u r   d u   a n v � n d e r ,   u n d e r h � l l e r   o c h   f e l s � k e r   d i n   p r o d u k t . "  
 F a s t F o t o   	 	 = " D e n   l � t e r   d i g   s n a b b t   s k a n n a   f o t o n   o c h   d o k u m e n t   o c h   � v e n   k o r r i g e r a   o c h   � t e r s t � l l a   f o t o n   s o m   � r   i   d � l i g t   s k i c k ,   s a m t   d e l a   d e m   e n k e l t . "  
 F a s t F o t o 2   	 	 = " D e n   l � t e r   d i g   s n a b b t   s k a n n a   f o t o n   o c h   d o k u m e n t   o c h   � v e n   k o r r i g e r a   o c h   � t e r s t � l l a   f o t o n   s o m   � r   i   d � l i g t   s k i c k ,   s a m t   d e l a   d e m   e n k e l t . "  
 S t a t u s M o n i t o r x 6 4 	 = " D e t   � v e r v a k a r   d i n   p r o d u k t   o c h   g e r   d i g   i n f o r m a t i o n   o m   s i n   s t a t u s . "  
 S t a t u s M o n i t o r x 8 6 	 = " D e t   � v e r v a k a r   d i n   p r o d u k t   o c h   g e r   d i g   i n f o r m a t i o n   o m   s i n   s t a t u s . "  
 S t a t u s M o n i t o r 3 	 	 = " D e t   � v e r v a k a r   d i n   p r o d u k t   o c h   g e r   d i g   i n f o r m a t i o n   o m   s i n   s t a t u s . "  
 C o n n e c t C h e c k e r   	 	 = " D e n   k o n t r o l l e r a r   s k r i v a r s t a t u s   o c h   f � r s � k e r   � t e r s t � l l a   u t s k r i f t   n � r   d e t   f i n n s   u t s k r i f t s p r o b l e m . "  
 P L o g A g e n t   	 	 = " D e t t a   � r   e t t   E p s o n   g l o b a l   r e s e a r c h - p r o g r a m   s o m   s a m l a r   i n   i n f o r m a t i o n   o m   d i n   p r o d u k t   s �   a t t   v i   k a n   f � r b � t t r a   v � r a   f r a m t i d a   p r o d u k t e r   o c h   t j � n s t e r .   V i   s a m l a r   i n t e   i n   p r o d u k t i n f o r m a t i o n   o m   d u   i n t e   g o d k � n n e r   d e t . "  
 S c a n S m a r t I J P   	 	 = " D e t   l � t e r   d i g   s k a n n a   d e t   u r s p r u n g l i g a   d o k u m e n t e t   o c h   s e d a n   f � l j a   i n s t r u k t i o n e r n a   p �   s k � r m e n   f � r   a t t   s p a r a   e l l e r   s k i c k a   d e n   s k a n n a d e   b i l d e n . "  
 D o c u m e n t C a p t u r e P r o V 2 I J P 	 = " D e t   l � t e r   d i g   h a n t e r a   s k a n n a d e   d o k u m e n t   o c h   s p a r a   d e m   s o m   f i l e r   f � r   a t t   s e d a n   s k i c k a   d e m   t i l l   F T P ,   e n   s k r i v a r e   e l l e r   m o l n e t . "  
 P r i n t e r D r i v e r x 6 4 _ L a b e l   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 P r i n t e r D r i v e r x 8 6 _ L a b e l   	 = " D e t   l � t e r   d i g   s t y r a   a l l a   a s p e k t e r   a v   u t s k r i f t ,   i n s t � l l n i n g a r   f � r   p a p p e r s t y p   o c h   p a p p e r s s t o r l e k ,   u t s k r i f t s k v a l i t e t   o c h   s �   v i d a r e . "  
 